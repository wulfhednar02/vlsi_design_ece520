* Circuit Extracted by Tanner Research's L-Edit V7.12 / Extract V4.00 ;
* TDB File:  C:\Users\ibows\Documents\ECE520\Project\Layout\Project_Inverter_v7, Cell:  Transceiver
* Extract Definition File:  ON_C5N.ext
* Extract Date and Time:  03/17/2019 - 23:53

.INCLUDE ON_C5N.modlib

* WARNING:  Layers with Unassigned AREA Capacitance.
*   <Substrate>
*   <ChipSubstrate>
* WARNING:  Layers with Unassigned FRINGE Capacitance.
*   <ndiff>
*   <Substrate>
*   <pdiff>
*   <n well wire>
*   <ChipSubstrate>
* WARNING:  Layers with Zero Resistance.
*   <Substrate>
*   <ChipSubstrate>

.subckt TRANSCEIVER TX RX CHANNEL VDD GND
* NODE NAME ALIASES
*       1 = GND (-241,-37.5)
*       1 = U10/GND (-19,-36.5)
*       1 = U11/GND (240,-38.5)
*       1 = U12/GND (269,-36)
*       1 = U16/GND (48,-36)
*       1 = U18/GND (296,-36)
*       1 = U23/GND (97,-36.5)
*       1 = U24/GND (213,-36)
*       1 = U35/GND (-241,-36)
*       1 = U36/GND (164,-36)
*       1 = U43/GND (-192,-36)
*       1 = U44/GND (-113,-36.5)
*       1 = U46/GND (-46,-36)
*       1 = U9/GND (-143,-36.5)
*       2 = VDD (-241,40.5)
*       2 = U10/VDD (-19,37.5)
*       2 = U11/VDD (240,39.5)
*       2 = U12/VDD (269,37)
*       2 = U16/VDD (48,37)
*       2 = U18/VDD (296,37)
*       2 = U23/VDD (97,37.5)
*       2 = U24/VDD (213,37)
*       2 = U35/VDD (-241,37)
*       2 = U36/VDD (164,37)
*       2 = U43/VDD (-192,37)
*       2 = U44/VDD (-113,37.5)
*       2 = U46/VDD (-46,37)
*       2 = U9/VDD (-143,37.5)
*       4 = CHANNEL (-241,56)
*       4 = U10/Input (-13.5,0.5)
*       4 = U43/Output (-147,0.5)
*       4 = U9/Input (-143,0.5)
*       5 = U23/Input (102.5,0.5)
*       5 = U35/Output (-196,0.5)
*       5 = U43/Input (-188,0.5)
*       7 = TX (-237,1)
*       7 = U35/Input (-237,0.5)
*       8 = U44/Input (-107.5,0.5)
*       8 = U9/Output (-119,0.5)
*       9 = U44/Output (-56,0.5)
*       9 = U46/Input (-42,0.5)
*       10 = U11/Select (243,0.5)
*       10 = U24/Output (236,0.5)
*       11 = U24/Input (217,0.5)
*       11 = U36/Output (209,0.5)
*       12 = U10/Output (38,0.5)
*       12 = U16/Input (52,0.5)
*       13 = U23/Output (154,0.5)
*       13 = U36/Input (168,0.5)
*       14 = U11/Input_N (243,-6)
*       14 = U16/Output (93,0.5)
*       17 = RX (340,1)
*       17 = U18/Output (341,0.5)
*       19 = U12/Output (292,0.5)
*       19 = U18/Input (300,0.5)
*       20 = U11/Output (263,0.5)
*       20 = U12/Input (273,0.5)
*       21 = U11/Input_P (243,7)
*       21 = U46/Output (-23,0.5)

Cpar1 GND 0 394.24689f
Cpar2 VDD 0 1.0803086p
Cpar3 3 0 27.073103f
Cpar4 CHANNEL 0 38.053287f
Cpar5 U23/Input 0 42.461476f
Cpar6 6 0 31.803217f
Cpar7 TX 0 1.0382228f
Cpar8 U44/Input 0 38.122681f
Cpar9 U44/Output 0 95.659303f
Cpar10 U11/Select 0 32.188599f
Cpar11 U24/Input 0 31.85453f
Cpar12 U10/Output 0 95.659303f
Cpar13 U23/Output 0 95.659303f
Cpar14 U11/Input_N 0 54.753238f
Cpar15 15 0 31.803217f
Cpar16 16 0 31.803217f
Cpar17 RX 0 30.744477f
Cpar18 18 0 31.803217f
Cpar19 U12/Output 0 31.85453f
Cpar20 U11/Output 0 60.141116f
Cpar21 U11/Input_P 0 56.020281f

M22 CHANNEL 3 VDD VDD CMOSP L=0.6u W=5.25u AD=8.6625p PD=13.8u AS=315.5625p PS=461.1u 
* M22 DRAIN GATE SOURCE BULK (-156.5 7.5 -154.5 25) 
M23 3 U23/Input VDD VDD CMOSP L=0.6u W=5.25u AD=8.6625p PD=13.8u AS=315.5625p PS=461.1u 
* M23 DRAIN GATE SOURCE BULK (-178.5 7.5 -176.5 25) 
M24 U23/Input 6 VDD VDD CMOSP L=0.6u W=6.75u AD=11.1375p PD=16.8u AS=315.5625p PS=461.1u 
* M24 DRAIN GATE SOURCE BULK (-205.5 6 -203.5 28.5) 
M25 6 TX VDD VDD CMOSP L=0.6u W=6.75u AD=11.1375p PD=16.8u AS=315.5625p PS=461.1u 
* M25 DRAIN GATE SOURCE BULK (-227.5 6 -225.5 28.5) 
M26 U44/Input CHANNEL VDD VDD CMOSP L=0.6u W=3u AD=4.95p PD=9.3u AS=315.5625p PS=461.1u 
* M26 DRAIN GATE SOURCE BULK (-129.5 6.5 -127.5 16.5) 
M27 VDD U44/Input U44/Output VDD CMOSP L=0.6u W=8.25u AD=315.5625p PD=461.1u AS=44.55p PS=60.3u 
* M27 DRAIN GATE SOURCE BULK (-59.5 6 -57.5 33.5) 
M28 U44/Output U44/Input VDD VDD CMOSP L=0.6u W=8.25u AD=44.55p PD=60.3u AS=315.5625p PS=461.1u 
* M28 DRAIN GATE SOURCE BULK (-67.5 6 -65.5 33.5) 
M29 VDD U44/Input U44/Output VDD CMOSP L=0.6u W=8.25u AD=315.5625p PD=461.1u AS=44.55p PS=60.3u 
* M29 DRAIN GATE SOURCE BULK (-75.5 6 -73.5 33.5) 
M30 U44/Output U44/Input VDD VDD CMOSP L=0.6u W=8.25u AD=44.55p PD=60.3u AS=315.5625p PS=461.1u 
* M30 DRAIN GATE SOURCE BULK (-83.5 6 -81.5 33.5) 
M31 VDD U44/Input U44/Output VDD CMOSP L=0.6u W=8.25u AD=315.5625p PD=461.1u AS=44.55p PS=60.3u 
* M31 DRAIN GATE SOURCE BULK (-91.5 6 -89.5 33.5) 
M32 U44/Output U44/Input VDD VDD CMOSP L=0.6u W=8.25u AD=44.55p PD=60.3u AS=315.5625p PS=461.1u 
* M32 DRAIN GATE SOURCE BULK (-99.5 6 -97.5 33.5) 
M33 U11/Input_P U44/Output VDD VDD CMOSP L=0.6u W=6.75u AD=22.5225p PD=33.9u AS=315.5625p PS=461.1u 
* M33 DRAIN GATE SOURCE BULK (-32.5 6 -30.5 28.5) 
M34 U11/Select U24/Input VDD VDD CMOSP L=0.6u W=6.75u AD=11.1375p PD=16.8u AS=315.5625p PS=461.1u 
* M34 DRAIN GATE SOURCE BULK (226.5 6 228.5 28.5) 
M35 VDD CHANNEL U10/Output VDD CMOSP L=0.6u W=8.25u AD=315.5625p PD=461.1u AS=44.55p PS=60.3u 
* M35 DRAIN GATE SOURCE BULK (34.5 6 36.5 33.5) 
M36 U10/Output CHANNEL VDD VDD CMOSP L=0.6u W=8.25u AD=44.55p PD=60.3u AS=315.5625p PS=461.1u 
* M36 DRAIN GATE SOURCE BULK (26.5 6 28.5 33.5) 
M37 VDD CHANNEL U10/Output VDD CMOSP L=0.6u W=8.25u AD=315.5625p PD=461.1u AS=44.55p PS=60.3u 
* M37 DRAIN GATE SOURCE BULK (18.5 6 20.5 33.5) 
M38 U10/Output CHANNEL VDD VDD CMOSP L=0.6u W=8.25u AD=44.55p PD=60.3u AS=315.5625p PS=461.1u 
* M38 DRAIN GATE SOURCE BULK (10.5 6 12.5 33.5) 
M39 VDD CHANNEL U10/Output VDD CMOSP L=0.6u W=8.25u AD=315.5625p PD=461.1u AS=44.55p PS=60.3u 
* M39 DRAIN GATE SOURCE BULK (2.5 6 4.5 33.5) 
M40 U10/Output CHANNEL VDD VDD CMOSP L=0.6u W=8.25u AD=44.55p PD=60.3u AS=315.5625p PS=461.1u 
* M40 DRAIN GATE SOURCE BULK (-5.5 6 -3.5 33.5) 
M41 VDD U23/Input U23/Output VDD CMOSP L=0.6u W=8.25u AD=315.5625p PD=461.1u AS=44.55p PS=60.3u 
* M41 DRAIN GATE SOURCE BULK (150.5 6 152.5 33.5) 
M42 U23/Output U23/Input VDD VDD CMOSP L=0.6u W=8.25u AD=44.55p PD=60.3u AS=315.5625p PS=461.1u 
* M42 DRAIN GATE SOURCE BULK (142.5 6 144.5 33.5) 
M43 VDD U23/Input U23/Output VDD CMOSP L=0.6u W=8.25u AD=315.5625p PD=461.1u AS=44.55p PS=60.3u 
* M43 DRAIN GATE SOURCE BULK (134.5 6 136.5 33.5) 
M44 U23/Output U23/Input VDD VDD CMOSP L=0.6u W=8.25u AD=44.55p PD=60.3u AS=315.5625p PS=461.1u 
* M44 DRAIN GATE SOURCE BULK (126.5 6 128.5 33.5) 
M45 VDD U23/Input U23/Output VDD CMOSP L=0.6u W=8.25u AD=315.5625p PD=461.1u AS=44.55p PS=60.3u 
* M45 DRAIN GATE SOURCE BULK (118.5 6 120.5 33.5) 
M46 U23/Output U23/Input VDD VDD CMOSP L=0.6u W=8.25u AD=44.55p PD=60.3u AS=315.5625p PS=461.1u 
* M46 DRAIN GATE SOURCE BULK (110.5 6 112.5 33.5) 
M47 U11/Input_N 15 VDD VDD CMOSP L=0.6u W=6.75u AD=11.1375p PD=16.8u AS=315.5625p PS=461.1u 
* M47 DRAIN GATE SOURCE BULK (83.5 6 85.5 28.5) 
M48 15 U10/Output VDD VDD CMOSP L=0.6u W=6.75u AD=11.1375p PD=16.8u AS=315.5625p PS=461.1u 
* M48 DRAIN GATE SOURCE BULK (61.5 6 63.5 28.5) 
M49 U24/Input 16 VDD VDD CMOSP L=0.6u W=6.75u AD=11.1375p PD=16.8u AS=315.5625p PS=461.1u 
* M49 DRAIN GATE SOURCE BULK (199.5 6 201.5 28.5) 
M50 16 U23/Output VDD VDD CMOSP L=0.6u W=6.75u AD=11.1375p PD=16.8u AS=315.5625p PS=461.1u 
* M50 DRAIN GATE SOURCE BULK (177.5 6 179.5 28.5) 
M51 RX 18 VDD VDD CMOSP L=0.6u W=6.75u AD=11.1375p PD=16.8u AS=315.5625p PS=461.1u 
* M51 DRAIN GATE SOURCE BULK (331.5 6 333.5 28.5) 
M52 18 U12/Output VDD VDD CMOSP L=0.6u W=6.75u AD=11.1375p PD=16.8u AS=315.5625p PS=461.1u 
* M52 DRAIN GATE SOURCE BULK (309.5 6 311.5 28.5) 
M53 U11/Output U11/Select U11/Input_P VDD CMOSP L=0.6u W=6.9u AD=15.525p PD=18.3u AS=22.5225p PS=33.9u 
* M53 DRAIN GATE SOURCE BULK (251.5 10.5 253.5 33.5) 
M54 U12/Output U11/Output VDD VDD CMOSP L=0.6u W=6.75u AD=11.1375p PD=16.8u AS=315.5625p PS=461.1u 
* M54 DRAIN GATE SOURCE BULK (282.5 6 284.5 28.5) 
M55 CHANNEL 3 GND GND CMOSN L=0.6u W=3u AD=4.95p PD=9.3u AS=99.99p PS=180.6u 
* M55 DRAIN GATE SOURCE BULK (-156.5 -17.5 -154.5 -7.5) 
M56 3 U23/Input GND GND CMOSN L=0.6u W=3u AD=4.95p PD=9.3u AS=99.99p PS=180.6u 
* M56 DRAIN GATE SOURCE BULK (-178.5 -17.5 -176.5 -7.5) 
M57 U23/Input 6 GND GND CMOSN L=0.6u W=3u AD=4.95p PD=9.3u AS=99.99p PS=180.6u 
* M57 DRAIN GATE SOURCE BULK (-205.5 -16 -203.5 -6) 
M58 6 TX GND GND CMOSN L=0.6u W=3u AD=4.95p PD=9.3u AS=99.99p PS=180.6u 
* M58 DRAIN GATE SOURCE BULK (-227.5 -16 -225.5 -6) 
M59 GND CHANNEL U44/Input GND CMOSN L=0.6u W=6.3u AD=99.99p PD=180.6u AS=11.34p PS=16.2u 
* M59 DRAIN GATE SOURCE BULK (-122.5 -27 -120.5 -6) 
M60 U44/Input CHANNEL GND GND CMOSN L=0.6u W=6.3u AD=11.34p PD=16.2u AS=99.99p PS=180.6u 
* M60 DRAIN GATE SOURCE BULK (-130.5 -27 -128.5 -6) 
M61 U44/Output U44/Input GND GND CMOSN L=3.6u W=3u AD=4.95p PD=9.3u AS=99.99p PS=180.6u 
* M61 DRAIN GATE SOURCE BULK (-77.5 -16.5 -65.5 -6.5) 
M62 U11/Input_P U44/Output GND GND CMOSN L=0.6u W=3u AD=4.95p PD=9.3u AS=99.99p PS=180.6u 
* M62 DRAIN GATE SOURCE BULK (-32.5 -16 -30.5 -6) 
M63 U11/Select U24/Input GND GND CMOSN L=0.6u W=3u AD=4.95p PD=9.3u AS=99.99p PS=180.6u 
* M63 DRAIN GATE SOURCE BULK (226.5 -16 228.5 -6) 
M64 U10/Output CHANNEL GND GND CMOSN L=3.6u W=3u AD=4.95p PD=9.3u AS=99.99p PS=180.6u 
* M64 DRAIN GATE SOURCE BULK (16.5 -16.5 28.5 -6.5) 
M65 U23/Output U23/Input GND GND CMOSN L=3.6u W=3u AD=4.95p PD=9.3u AS=99.99p PS=180.6u 
* M65 DRAIN GATE SOURCE BULK (132.5 -16.5 144.5 -6.5) 
M66 U11/Input_N 15 GND GND CMOSN L=0.6u W=3u AD=16.335p PD=26.4u AS=99.99p PS=180.6u 
* M66 DRAIN GATE SOURCE BULK (83.5 -16 85.5 -6) 
M67 15 U10/Output GND GND CMOSN L=0.6u W=3u AD=4.95p PD=9.3u AS=99.99p PS=180.6u 
* M67 DRAIN GATE SOURCE BULK (61.5 -16 63.5 -6) 
M68 U24/Input 16 GND GND CMOSN L=0.6u W=3u AD=4.95p PD=9.3u AS=99.99p PS=180.6u 
* M68 DRAIN GATE SOURCE BULK (199.5 -16 201.5 -6) 
M69 16 U23/Output GND GND CMOSN L=0.6u W=3u AD=4.95p PD=9.3u AS=99.99p PS=180.6u 
* M69 DRAIN GATE SOURCE BULK (177.5 -16 179.5 -6) 
M70 RX 18 GND GND CMOSN L=0.6u W=3u AD=4.95p PD=9.3u AS=99.99p PS=180.6u 
* M70 DRAIN GATE SOURCE BULK (331.5 -16 333.5 -6) 
M71 18 U12/Output GND GND CMOSN L=0.6u W=3u AD=4.95p PD=9.3u AS=99.99p PS=180.6u 
* M71 DRAIN GATE SOURCE BULK (309.5 -16 311.5 -6) 
M72 U11/Output U11/Select U11/Input_N GND CMOSN L=0.6u W=6.9u AD=15.525p PD=18.3u AS=16.335p PS=26.4u 
* M72 DRAIN GATE SOURCE BULK (251.5 -33.5 253.5 -10.5) 
M73 U12/Output U11/Output GND GND CMOSN L=0.6u W=3u AD=4.95p PD=9.3u AS=99.99p PS=180.6u 
* M73 DRAIN GATE SOURCE BULK (282.5 -16 284.5 -6) 
.ends

Vsupply VDD 0 5

* transceiver 1
Xtrans1 TX1 RX1 channel VDD 0 TRANSCEIVER
* transceiver 2
Xtrans2 TX2 RX2 channel VDD 0 TRANSCEIVER

* pad, etc. loads on receiver output
*Crx1load RX1 0 20p
*Crx2load RX2 0 20p

* Input waveforms as stimulus
Vtx1 TX1 0 PULSE(0 5 0 10n 10n 100n 400n)
Vtx2 TX2 0 PULSE(0 5 0 10n 10n 30n 90n)

.probe

.tran 1p 2u

* Total Nodes: 21
* Total Elements: 73
* Extract Elapsed Time: 0 seconds
.END
