.SUBCKT 2TMUX P_IN N_IN SEL OUT VDD GND

* if (sel==0) out=P_IN
* else out=N_IN

Mp OUT SEL P_IN VDD CMOSP L=0.6u W={MIN_CHANNEL_WIDTH*BALANCED_RATIO} PS=8.4u PD=8.4u
Mn OUT SEL N_IN GND CMOSN L=0.6u W={MIN_CHANNEL_WIDTH} PS=8.4u PD=8.4u
.ENDS
