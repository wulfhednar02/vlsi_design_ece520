
.SUBCKT INVX9 IN OUT VDD GND

* NODE NAME ALIASES
*       1 = GND (49.499,-56.499)
*       2 = VDD (-46.5,77.5)
*       3 = INVX1 (-24,17.5)
*       4 = OUT (63.499,-7.999)
*       5 = INVX3 (0,19.5)
*       6 = IN (-35,17)

Cpar1 GND 0 273.33037f
Cpar2 VDD 0 423.23035f
Cpar3 INVX1 0 39.20328f
Cpar4 OUT 0 302.38707f
Cpar5 INVX3 0 112.49626f
Cpar6 IN 0 5.0056642f
Cpar7 7 0 53.7075f

M8 OUT INVX3 VDD 7 CMOSP L=0.6u W=14.85u AD=98.01p PD=72.6u AS=218.3175p PS=171.3u 
* M8 DRAIN GATE SOURCE BULK (54.5 14.5 56.5 64) 
M9 OUT INVX3 VDD 7 CMOSP L=0.6u W=14.85u AD=98.01p PD=72.6u AS=218.3175p PS=171.3u 
* M9 DRAIN GATE SOURCE BULK (41.5 14.5 43.5 64) 
M10 OUT INVX3 VDD 7 CMOSP L=0.6u W=14.85u AD=98.01p PD=72.6u AS=218.3175p PS=171.3u 
* M10 DRAIN GATE SOURCE BULK (28.5 14.5 30.5 64) 
M11 OUT INVX3 VDD 7 CMOSP L=0.6u W=14.85u AD=98.01p PD=72.6u AS=218.3175p PS=171.3u 
* M11 DRAIN GATE SOURCE BULK (15.5 14.5 17.5 64) 
M12 INVX3 INVX1 VDD 7 CMOSP L=0.6u W=9.9u AD=32.67p PD=26.4u AS=218.3175p PS=171.3u 
* M12 DRAIN GATE SOURCE BULK (-2.5 31 -0.5 64) 
M13 INVX3 INVX1 VDD 7 CMOSP L=0.6u W=9.9u AD=32.67p PD=26.4u AS=218.3175p PS=171.3u 
* M13 DRAIN GATE SOURCE BULK (-15.5 31 -13.5 64) 
M14 INVX1 IN VDD 7 CMOSP L=0.6u W=3.3u AD=5.94p PD=10.2u AS=218.3175p PS=171.3u 
* M14 DRAIN GATE SOURCE BULK (-31.5 53 -29.5 64) 
M15 INVX1 IN VDD 7 CMOSP L=0.6u W=3.3u AD=5.94p PD=10.2u AS=218.3175p PS=171.3u 
* M15 DRAIN GATE SOURCE BULK (-39.5 53 -37.5 64) 
M16 OUT INVX3 GND GND CMOSN L=0.6u W=9u AD=59.4p PD=49.2u AS=99.135p PS=94.8u 
* M16 DRAIN GATE SOURCE BULK (45.5 -46 47.5 -16) 
M17 OUT INVX3 GND GND CMOSN L=0.6u W=9u AD=59.4p PD=49.2u AS=99.135p PS=94.8u 
* M17 DRAIN GATE SOURCE BULK (32.5 -46 34.5 -16) 
M18 OUT INVX3 GND GND CMOSN L=0.6u W=9u AD=59.4p PD=49.2u AS=99.135p PS=94.8u 
* M18 DRAIN GATE SOURCE BULK (19.5 -46 21.5 -16) 
M19 INVX3 INVX1 GND GND CMOSN L=0.6u W=4.5u AD=16.2p PD=16.2u AS=99.135p PS=94.8u 
* M19 DRAIN GATE SOURCE BULK (6 -40.5 8 -25.5) 
M20 INVX3 INVX1 GND GND CMOSN L=0.6u W=4.5u AD=16.2p PD=16.2u AS=99.135p PS=94.8u 
* M20 DRAIN GATE SOURCE BULK (-8 -40.5 -6 -25.5) 
M21 INVX1 IN GND GND CMOSN L=0.6u W=3u AD=10.35p PD=12.9u AS=99.135p PS=94.8u 
* M21 DRAIN GATE SOURCE BULK (-37 -36 -35 -26) 

* Total Nodes: 7
* Total Elements: 21
* Extract Elapsed Time: 0 seconds

.ENDS
