.SUBCKT 2TMUX P_IN N_IN SEL OUT VDD GND

* if (sel==0) out=P_IN
* else out=N_IN

Mp OUT SEL P_IN VDD CMOSP 
+L=0.6u 
+W={MIN_CHANNEL_WIDTH*BALANCED_RATIO} 
+AS=(BALANCED_RATIO*MIN_CHANNEL_WIDTH*1.5u)
+AD=(BALANCED_RATIO*MIN_CHANNEL_WIDTH*1.5u)
+PS=(8.4u+((BALANCED_RATIO-1)*MIN_CHANNEL_WIDTH))
+PD=(8.4u+((BALANCED_RATIO-1)*MIN_CHANNEL_WIDTH))

Mn OUT SEL N_IN GND CMOSN
+L=0.6u
+W={MIN_CHANNEL_WIDTH}
+AS=4.5p
+AD=4.5p
+PS=8.4u
+PD=8.4u

.ENDS
