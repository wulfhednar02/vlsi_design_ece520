
.SUBCKT INVX81 IN OUT VDD GND

* NODE NAME ALIASES
*       1 = GND (58.667,148)
*       2 = VDD (4.667,7)
*       3 = IN (341.666,99)
*       4 = OUT (38.666,96)

Cpar1 GND 0 1.5499151p
Cpar2 VDD 0 2.4134859p
Cpar3 IN 0 84.693252f
Cpar4 OUT 0 2.4832353p

M5 OUT IN VDD VDD CMOSP L=0.6u W=22.35u AD=885.06p PD=615.6u AS=996.9525p PS=691.2u 
* M5 DRAIN GATE SOURCE BULK (321.667 14 323.667 88.5) 
M6 OUT IN VDD VDD CMOSP L=0.6u W=22.35u AD=885.06p PD=615.6u AS=996.9525p PS=691.2u 
* M6 DRAIN GATE SOURCE BULK (308.667 14 310.667 88.5) 
M7 OUT IN VDD VDD CMOSP L=0.6u W=22.35u AD=885.06p PD=615.6u AS=996.9525p PS=691.2u 
* M7 DRAIN GATE SOURCE BULK (295.667 14 297.667 88.5) 
M8 OUT IN VDD VDD CMOSP L=0.6u W=22.35u AD=885.06p PD=615.6u AS=996.9525p PS=691.2u 
* M8 DRAIN GATE SOURCE BULK (282.667 14 284.667 88.5) 
M9 OUT IN VDD VDD CMOSP L=0.6u W=22.35u AD=885.06p PD=615.6u AS=996.9525p PS=691.2u 
* M9 DRAIN GATE SOURCE BULK (269.667 14 271.667 88.5) 
M10 OUT IN VDD VDD CMOSP L=0.6u W=22.35u AD=885.06p PD=615.6u AS=996.9525p PS=691.2u 
* M10 DRAIN GATE SOURCE BULK (256.667 14 258.667 88.5) 
M11 OUT IN VDD VDD CMOSP L=0.6u W=22.35u AD=885.06p PD=615.6u AS=996.9525p PS=691.2u 
* M11 DRAIN GATE SOURCE BULK (243.667 14 245.667 88.5) 
M12 OUT IN VDD VDD CMOSP L=0.6u W=22.35u AD=885.06p PD=615.6u AS=996.9525p PS=691.2u 
* M12 DRAIN GATE SOURCE BULK (230.667 14 232.667 88.5) 
M13 OUT IN VDD VDD CMOSP L=0.6u W=22.35u AD=885.06p PD=615.6u AS=996.9525p PS=691.2u 
* M13 DRAIN GATE SOURCE BULK (217.667 14 219.667 88.5) 
M14 OUT IN VDD VDD CMOSP L=0.6u W=22.35u AD=885.06p PD=615.6u AS=996.9525p PS=691.2u 
* M14 DRAIN GATE SOURCE BULK (204.667 14 206.667 88.5) 
M15 OUT IN VDD VDD CMOSP L=0.6u W=22.35u AD=885.06p PD=615.6u AS=996.9525p PS=691.2u 
* M15 DRAIN GATE SOURCE BULK (191.667 14 193.667 88.5) 
M16 OUT IN VDD VDD CMOSP L=0.6u W=22.35u AD=885.06p PD=615.6u AS=996.9525p PS=691.2u 
* M16 DRAIN GATE SOURCE BULK (178.667 14 180.667 88.5) 
M17 OUT IN VDD VDD CMOSP L=0.6u W=22.35u AD=885.06p PD=615.6u AS=996.9525p PS=691.2u 
* M17 DRAIN GATE SOURCE BULK (165.667 14 167.667 88.5) 
M18 OUT IN VDD VDD CMOSP L=0.6u W=22.35u AD=885.06p PD=615.6u AS=996.9525p PS=691.2u 
* M18 DRAIN GATE SOURCE BULK (152.667 14 154.667 88.5) 
M19 OUT IN VDD VDD CMOSP L=0.6u W=22.35u AD=885.06p PD=615.6u AS=996.9525p PS=691.2u 
* M19 DRAIN GATE SOURCE BULK (139.667 14 141.667 88.5) 
M20 OUT IN VDD VDD CMOSP L=0.6u W=22.35u AD=885.06p PD=615.6u AS=996.9525p PS=691.2u 
* M20 DRAIN GATE SOURCE BULK (126.667 14 128.667 88.5) 
M21 OUT IN VDD VDD CMOSP L=0.6u W=22.35u AD=885.06p PD=615.6u AS=996.9525p PS=691.2u 
* M21 DRAIN GATE SOURCE BULK (113.667 14 115.667 88.5) 
M22 OUT IN VDD VDD CMOSP L=0.6u W=22.35u AD=885.06p PD=615.6u AS=996.9525p PS=691.2u 
* M22 DRAIN GATE SOURCE BULK (100.667 14 102.667 88.5) 
M23 OUT IN VDD VDD CMOSP L=0.6u W=22.35u AD=885.06p PD=615.6u AS=996.9525p PS=691.2u 
* M23 DRAIN GATE SOURCE BULK (87.667 14 89.667 88.5) 
M24 OUT IN VDD VDD CMOSP L=0.6u W=22.35u AD=885.06p PD=615.6u AS=996.9525p PS=691.2u 
* M24 DRAIN GATE SOURCE BULK (74.667 14 76.667 88.5) 
M25 OUT IN VDD VDD CMOSP L=0.6u W=22.35u AD=885.06p PD=615.6u AS=996.9525p PS=691.2u 
* M25 DRAIN GATE SOURCE BULK (61.667 14 63.667 88.5) 
M26 OUT IN VDD VDD CMOSP L=0.6u W=22.35u AD=885.06p PD=615.6u AS=996.9525p PS=691.2u 
* M26 DRAIN GATE SOURCE BULK (48.667 14 50.667 88.5) 
M27 OUT IN VDD VDD CMOSP L=0.6u W=22.35u AD=885.06p PD=615.6u AS=996.9525p PS=691.2u 
* M27 DRAIN GATE SOURCE BULK (35.667 14 37.667 88.5) 
M28 OUT IN VDD VDD CMOSP L=0.6u W=22.35u AD=885.06p PD=615.6u AS=996.9525p PS=691.2u 
* M28 DRAIN GATE SOURCE BULK (22.667 14 24.667 88.5) 
M29 OUT IN GND GND CMOSN L=0.6u W=10.2u AD=403.92p PD=324u AS=464.13p PS=374.1u 
* M29 DRAIN GATE SOURCE BULK (321.667 104.5 323.667 138.5) 
M30 OUT IN GND GND CMOSN L=0.6u W=10.2u AD=403.92p PD=324u AS=464.13p PS=374.1u 
* M30 DRAIN GATE SOURCE BULK (308.667 104.5 310.667 138.5) 
M31 OUT IN GND GND CMOSN L=0.6u W=10.2u AD=403.92p PD=324u AS=464.13p PS=374.1u 
* M31 DRAIN GATE SOURCE BULK (295.667 104.5 297.667 138.5) 
M32 OUT IN GND GND CMOSN L=0.6u W=10.2u AD=403.92p PD=324u AS=464.13p PS=374.1u 
* M32 DRAIN GATE SOURCE BULK (282.667 104.5 284.667 138.5) 
M33 OUT IN GND GND CMOSN L=0.6u W=10.2u AD=403.92p PD=324u AS=464.13p PS=374.1u 
* M33 DRAIN GATE SOURCE BULK (269.667 104.5 271.667 138.5) 
M34 OUT IN GND GND CMOSN L=0.6u W=10.2u AD=403.92p PD=324u AS=464.13p PS=374.1u 
* M34 DRAIN GATE SOURCE BULK (256.667 104.5 258.667 138.5) 
M35 OUT IN GND GND CMOSN L=0.6u W=10.2u AD=403.92p PD=324u AS=464.13p PS=374.1u 
* M35 DRAIN GATE SOURCE BULK (243.667 104.5 245.667 138.5) 
M36 OUT IN GND GND CMOSN L=0.6u W=10.2u AD=403.92p PD=324u AS=464.13p PS=374.1u 
* M36 DRAIN GATE SOURCE BULK (230.667 104.5 232.667 138.5) 
M37 OUT IN GND GND CMOSN L=0.6u W=10.2u AD=403.92p PD=324u AS=464.13p PS=374.1u 
* M37 DRAIN GATE SOURCE BULK (217.667 104.5 219.667 138.5) 
M38 OUT IN GND GND CMOSN L=0.6u W=10.2u AD=403.92p PD=324u AS=464.13p PS=374.1u 
* M38 DRAIN GATE SOURCE BULK (204.667 104.5 206.667 138.5) 
M39 OUT IN GND GND CMOSN L=0.6u W=10.2u AD=403.92p PD=324u AS=464.13p PS=374.1u 
* M39 DRAIN GATE SOURCE BULK (191.667 104.5 193.667 138.5) 
M40 OUT IN GND GND CMOSN L=0.6u W=10.2u AD=403.92p PD=324u AS=464.13p PS=374.1u 
* M40 DRAIN GATE SOURCE BULK (178.667 104.5 180.667 138.5) 
M41 OUT IN GND GND CMOSN L=0.6u W=10.2u AD=403.92p PD=324u AS=464.13p PS=374.1u 
* M41 DRAIN GATE SOURCE BULK (165.667 104.5 167.667 138.5) 
M42 OUT IN GND GND CMOSN L=0.6u W=10.2u AD=403.92p PD=324u AS=464.13p PS=374.1u 
* M42 DRAIN GATE SOURCE BULK (152.667 104.5 154.667 138.5) 
M43 OUT IN GND GND CMOSN L=0.6u W=10.2u AD=403.92p PD=324u AS=464.13p PS=374.1u 
* M43 DRAIN GATE SOURCE BULK (139.667 104.5 141.667 138.5) 
M44 OUT IN GND GND CMOSN L=0.6u W=10.2u AD=403.92p PD=324u AS=464.13p PS=374.1u 
* M44 DRAIN GATE SOURCE BULK (126.667 104.5 128.667 138.5) 
M45 OUT IN GND GND CMOSN L=0.6u W=10.2u AD=403.92p PD=324u AS=464.13p PS=374.1u 
* M45 DRAIN GATE SOURCE BULK (113.667 104.5 115.667 138.5) 
M46 OUT IN GND GND CMOSN L=0.6u W=10.2u AD=403.92p PD=324u AS=464.13p PS=374.1u 
* M46 DRAIN GATE SOURCE BULK (100.667 104.5 102.667 138.5) 
M47 OUT IN GND GND CMOSN L=0.6u W=10.2u AD=403.92p PD=324u AS=464.13p PS=374.1u 
* M47 DRAIN GATE SOURCE BULK (87.667 104.5 89.667 138.5) 
M48 OUT IN GND GND CMOSN L=0.6u W=10.2u AD=403.92p PD=324u AS=464.13p PS=374.1u 
* M48 DRAIN GATE SOURCE BULK (74.667 104.5 76.667 138.5) 
M49 OUT IN GND GND CMOSN L=0.6u W=10.2u AD=403.92p PD=324u AS=464.13p PS=374.1u 
* M49 DRAIN GATE SOURCE BULK (61.667 104.5 63.667 138.5) 
M50 OUT IN GND GND CMOSN L=0.6u W=10.2u AD=403.92p PD=324u AS=464.13p PS=374.1u 
* M50 DRAIN GATE SOURCE BULK (48.667 104.5 50.667 138.5) 
M51 OUT IN GND GND CMOSN L=0.6u W=10.2u AD=403.92p PD=324u AS=464.13p PS=374.1u 
* M51 DRAIN GATE SOURCE BULK (35.667 104.5 37.667 138.5) 
M52 OUT IN GND GND CMOSN L=0.6u W=10.2u AD=403.92p PD=324u AS=464.13p PS=374.1u 
* M52 DRAIN GATE SOURCE BULK (22.667 104.5 24.667 138.5) 

.ENDS
