.SUBCKT INV_P_STRONG IN OUT VDD GND
.param X=1 * X is drive strength(width multiplier), as in INVX1, INVX4, etc.

* Vm = 3.75
* OUT = ~IN

Mp OUT IN VDD VDD CMOSP 
+L=0.6u
+W={X*MIN_CHANNEL_WIDTH*P_STRONG_RATIO}
+AS=(X*P_STRONG_RATIO*MIN_CHANNEL_WIDTH*1.5u)
+AD=(X*P_STRONG_RATIO*MIN_CHANNEL_WIDTH*1.5u)
+PS=(8.4u+(((X*P_STRONG_RATIO)-1)*MIN_CHANNEL_WIDTH))
+PD=(8.4u+(((X*P_STRONG_RATIO)-1)*MIN_CHANNEL_WIDTH))

Mn OUT IN GND GND CMOSN
+L=0.6u
+W={X*MIN_CHANNEL_WIDTH}
+AS=(X*MIN_CHANNEL_WIDTH*1.5u)
+AD=(X*MIN_CHANNEL_WIDTH*1.5u)
+PS=(8.4u+((X-1)*MIN_CHANNEL_WIDTH))
+PD=(8.4u+((X-1)*MIN_CHANNEL_WIDTH))

.ENDS
