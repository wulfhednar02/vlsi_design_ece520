
.INCLUDE INVX9.sp
.INCLUDE INVX27.sp
.INCLUDE INVX81.sp

.SUBCKT OUTBUF IN OUT VDD GND

Xinvx9 IN OUTX9 VDD GND INVX9
Xinvx27 OUTX9 OUTX27 VDD GND INVX27
Xinvx81 OUTX27 OUT VDD GND INVX81

.ENDS
