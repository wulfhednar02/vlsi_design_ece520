.SUBCKT INV_N_STRONG IN OUT VDD GND

* Vm = 3.75
* OUT = ~IN

Mp OUT IN VDD VDD CMOSP
+L=0.6u
+W={MIN_CHANNEL_WIDTH}
+AS=4.5p
+AD=4.5p
+PS=8.4u
+PD=8.4u

Mn OUT IN GND GND CMOSN
+L=0.6u
+W={MIN_CHANNEL_WIDTH*N_STRONG_RATIO}
+AS={N_STRONG_RATIO*MIN_CHANNEL_WIDTH*1.5u}
+AD={N_STRONG_RATIO*MIN_CHANNEL_WIDTH*1.5u}
+PS={8.4u+(((N_STRONG_RATIO)-1)*MIN_CHANNEL_WIDTH)}
+PD={8.4u+(((N_STRONG_RATIO)-1)*MIN_CHANNEL_WIDTH)}

.ENDS
