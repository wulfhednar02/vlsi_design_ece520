
.SUBCKT INVX27 IN OUT VDD GND

* WARNING: Node 1 has zero nodal parasitic capacitance.
Cpar1 GND 0 1.2799989p
Cpar2 VDD 0 669.62408f
Cpar3 IN 0 49.351431f
Cpar4 5 0 77.12397f

M5 VDD IN GND 5 CMOSP L=0.6u W=14.85u AD=345.2625p PD=254.4u AS=294.03p PS=217.8u 
* M5 DRAIN GATE SOURCE BULK (151.5 14.5 153.5 64) 
M6 GND IN VDD 5 CMOSP L=0.6u W=14.85u AD=294.03p PD=217.8u AS=345.2625p PS=254.4u 
* M6 DRAIN GATE SOURCE BULK (138.5 14.5 140.5 64) 
M7 VDD IN GND 5 CMOSP L=0.6u W=14.85u AD=345.2625p PD=254.4u AS=294.03p PS=217.8u 
* M7 DRAIN GATE SOURCE BULK (125.5 14.5 127.5 64) 
M8 GND IN VDD 5 CMOSP L=0.6u W=14.85u AD=294.03p PD=217.8u AS=345.2625p PS=254.4u 
* M8 DRAIN GATE SOURCE BULK (112.5 14.5 114.5 64) 
M9 VDD IN GND 5 CMOSP L=0.6u W=14.85u AD=345.2625p PD=254.4u AS=294.03p PS=217.8u 
* M9 DRAIN GATE SOURCE BULK (99 14.5 101 64) 
M10 GND IN VDD 5 CMOSP L=0.6u W=14.85u AD=294.03p PD=217.8u AS=345.2625p PS=254.4u 
* M10 DRAIN GATE SOURCE BULK (86 14.5 88 64) 
M11 VDD IN GND 5 CMOSP L=0.6u W=14.85u AD=345.2625p PD=254.4u AS=294.03p PS=217.8u 
* M11 DRAIN GATE SOURCE BULK (73 14.5 75 64) 
M12 GND IN VDD 5 CMOSP L=0.6u W=14.85u AD=294.03p PD=217.8u AS=345.2625p PS=254.4u 
* M12 DRAIN GATE SOURCE BULK (60 14.5 62 64) 
M13 VDD IN GND 5 CMOSP L=0.6u W=14.85u AD=345.2625p PD=254.4u AS=294.03p PS=217.8u 
* M13 DRAIN GATE SOURCE BULK (47 14.5 49 64) 
M14 GND IN VDD 5 CMOSP L=0.6u W=14.85u AD=294.03p PD=217.8u AS=345.2625p PS=254.4u 
* M14 DRAIN GATE SOURCE BULK (34 14.5 36 64) 
M15 VDD IN GND 5 CMOSP L=0.6u W=14.85u AD=345.2625p PD=254.4u AS=294.03p PS=217.8u 
* M15 DRAIN GATE SOURCE BULK (21 14.5 23 64) 
M16 GND IN VDD 5 CMOSP L=0.6u W=14.85u AD=294.03p PD=217.8u AS=345.2625p PS=254.4u 
* M16 DRAIN GATE SOURCE BULK (8 14.5 10 64) 
M17 GND IN GND 1 CMOSN L=0.6u W=9u AD=365.85p PD=261.3u AS=365.85p PS=261.3u 
* M17 DRAIN GATE SOURCE BULK (148.5 -46 150.5 -16) 
M18 GND IN GND 1 CMOSN L=0.6u W=9u AD=365.85p PD=261.3u AS=365.85p PS=261.3u 
* M18 DRAIN GATE SOURCE BULK (135.5 -46 137.5 -16) 
M19 GND IN GND 1 CMOSN L=0.6u W=9u AD=365.85p PD=261.3u AS=365.85p PS=261.3u 
* M19 DRAIN GATE SOURCE BULK (122.5 -46 124.5 -16) 
M20 GND IN GND 1 CMOSN L=0.6u W=9u AD=365.85p PD=261.3u AS=365.85p PS=261.3u 
* M20 DRAIN GATE SOURCE BULK (97 -46 99 -16) 
M21 GND IN GND 1 CMOSN L=0.6u W=9u AD=365.85p PD=261.3u AS=365.85p PS=261.3u 
* M21 DRAIN GATE SOURCE BULK (84 -46 86 -16) 
M22 GND IN GND 1 CMOSN L=0.6u W=9u AD=365.85p PD=261.3u AS=365.85p PS=261.3u 
* M22 DRAIN GATE SOURCE BULK (71 -46 73 -16) 
M23 GND IN GND 1 CMOSN L=0.6u W=9u AD=365.85p PD=261.3u AS=365.85p PS=261.3u 
* M23 DRAIN GATE SOURCE BULK (45.5 -46 47.5 -16) 
M24 GND IN GND 1 CMOSN L=0.6u W=9u AD=365.85p PD=261.3u AS=365.85p PS=261.3u 
* M24 DRAIN GATE SOURCE BULK (32.5 -46 34.5 -16) 
M25 GND IN GND 1 CMOSN L=0.6u W=9u AD=365.85p PD=261.3u AS=365.85p PS=261.3u 
* M25 DRAIN GATE SOURCE BULK (19.5 -46 21.5 -16) 

* Total Nodes: 5
* Total Elements: 25
* Extract Elapsed Time: 0 seconds
.ENDS
