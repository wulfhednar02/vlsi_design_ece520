
.SUBCKT INVX81 IN OUT VDD GND
Cpar1 GND 0 1.1727431p
Cpar2 VDD 0 2.369203p
Cpar3 IN 0 84.600904f
Cpar4 OUT 0 2.4832353p

M5 OUT IN GND GND CMOSN L=0.6u W=10.2u AD=403.92p PD=324u AS=464.13p PS=374.1u 
* M5 DRAIN GATE SOURCE BULK (322 104.5 324 138.5) 
M6 OUT IN GND GND CMOSN L=0.6u W=10.2u AD=403.92p PD=324u AS=464.13p PS=374.1u 
* M6 DRAIN GATE SOURCE BULK (309 104.5 311 138.5) 
M7 OUT IN GND GND CMOSN L=0.6u W=10.2u AD=403.92p PD=324u AS=464.13p PS=374.1u 
* M7 DRAIN GATE SOURCE BULK (296 104.5 298 138.5) 
M8 OUT IN GND GND CMOSN L=0.6u W=10.2u AD=403.92p PD=324u AS=464.13p PS=374.1u 
* M8 DRAIN GATE SOURCE BULK (283 104.5 285 138.5) 
M9 OUT IN GND GND CMOSN L=0.6u W=10.2u AD=403.92p PD=324u AS=464.13p PS=374.1u 
* M9 DRAIN GATE SOURCE BULK (270 104.5 272 138.5) 
M10 OUT IN GND GND CMOSN L=0.6u W=10.2u AD=403.92p PD=324u AS=464.13p PS=374.1u 
* M10 DRAIN GATE SOURCE BULK (257 104.5 259 138.5) 
M11 OUT IN GND GND CMOSN L=0.6u W=10.2u AD=403.92p PD=324u AS=464.13p PS=374.1u 
* M11 DRAIN GATE SOURCE BULK (244 104.5 246 138.5) 
M12 OUT IN GND GND CMOSN L=0.6u W=10.2u AD=403.92p PD=324u AS=464.13p PS=374.1u 
* M12 DRAIN GATE SOURCE BULK (231 104.5 233 138.5) 
M13 OUT IN GND GND CMOSN L=0.6u W=10.2u AD=403.92p PD=324u AS=464.13p PS=374.1u 
* M13 DRAIN GATE SOURCE BULK (218 104.5 220 138.5) 
M14 OUT IN GND GND CMOSN L=0.6u W=10.2u AD=403.92p PD=324u AS=464.13p PS=374.1u 
* M14 DRAIN GATE SOURCE BULK (205 104.5 207 138.5) 
M15 OUT IN GND GND CMOSN L=0.6u W=10.2u AD=403.92p PD=324u AS=464.13p PS=374.1u 
* M15 DRAIN GATE SOURCE BULK (192 104.5 194 138.5) 
M16 OUT IN GND GND CMOSN L=0.6u W=10.2u AD=403.92p PD=324u AS=464.13p PS=374.1u 
* M16 DRAIN GATE SOURCE BULK (179 104.5 181 138.5) 
M17 OUT IN GND GND CMOSN L=0.6u W=10.2u AD=403.92p PD=324u AS=464.13p PS=374.1u 
* M17 DRAIN GATE SOURCE BULK (166 104.5 168 138.5) 
M18 OUT IN GND GND CMOSN L=0.6u W=10.2u AD=403.92p PD=324u AS=464.13p PS=374.1u 
* M18 DRAIN GATE SOURCE BULK (153 104.5 155 138.5) 
M19 OUT IN GND GND CMOSN L=0.6u W=10.2u AD=403.92p PD=324u AS=464.13p PS=374.1u 
* M19 DRAIN GATE SOURCE BULK (140 104.5 142 138.5) 
M20 OUT IN GND GND CMOSN L=0.6u W=10.2u AD=403.92p PD=324u AS=464.13p PS=374.1u 
* M20 DRAIN GATE SOURCE BULK (127 104.5 129 138.5) 
M21 OUT IN GND GND CMOSN L=0.6u W=10.2u AD=403.92p PD=324u AS=464.13p PS=374.1u 
* M21 DRAIN GATE SOURCE BULK (114 104.5 116 138.5) 
M22 OUT IN GND GND CMOSN L=0.6u W=10.2u AD=403.92p PD=324u AS=464.13p PS=374.1u 
* M22 DRAIN GATE SOURCE BULK (101 104.5 103 138.5) 
M23 OUT IN GND GND CMOSN L=0.6u W=10.2u AD=403.92p PD=324u AS=464.13p PS=374.1u 
* M23 DRAIN GATE SOURCE BULK (88 104.5 90 138.5) 
M24 OUT IN GND GND CMOSN L=0.6u W=10.2u AD=403.92p PD=324u AS=464.13p PS=374.1u 
* M24 DRAIN GATE SOURCE BULK (75 104.5 77 138.5) 
M25 OUT IN GND GND CMOSN L=0.6u W=10.2u AD=403.92p PD=324u AS=464.13p PS=374.1u 
* M25 DRAIN GATE SOURCE BULK (62 104.5 64 138.5) 
M26 OUT IN GND GND CMOSN L=0.6u W=10.2u AD=403.92p PD=324u AS=464.13p PS=374.1u 
* M26 DRAIN GATE SOURCE BULK (49 104.5 51 138.5) 
M27 OUT IN GND GND CMOSN L=0.6u W=10.2u AD=403.92p PD=324u AS=464.13p PS=374.1u 
* M27 DRAIN GATE SOURCE BULK (36 104.5 38 138.5) 
M28 OUT IN GND GND CMOSN L=0.6u W=10.2u AD=403.92p PD=324u AS=464.13p PS=374.1u 
* M28 DRAIN GATE SOURCE BULK (23 104.5 25 138.5) 
M29 OUT IN VDD VDD CMOSP L=0.6u W=22.35u AD=885.06p PD=615.6u AS=996.9525p PS=691.2u 
* M29 DRAIN GATE SOURCE BULK (322 14 324 88.5) 
M30 OUT IN VDD VDD CMOSP L=0.6u W=22.35u AD=885.06p PD=615.6u AS=996.9525p PS=691.2u 
* M30 DRAIN GATE SOURCE BULK (309 14 311 88.5) 
M31 OUT IN VDD VDD CMOSP L=0.6u W=22.35u AD=885.06p PD=615.6u AS=996.9525p PS=691.2u 
* M31 DRAIN GATE SOURCE BULK (296 14 298 88.5) 
M32 OUT IN VDD VDD CMOSP L=0.6u W=22.35u AD=885.06p PD=615.6u AS=996.9525p PS=691.2u 
* M32 DRAIN GATE SOURCE BULK (283 14 285 88.5) 
M33 OUT IN VDD VDD CMOSP L=0.6u W=22.35u AD=885.06p PD=615.6u AS=996.9525p PS=691.2u 
* M33 DRAIN GATE SOURCE BULK (270 14 272 88.5) 
M34 OUT IN VDD VDD CMOSP L=0.6u W=22.35u AD=885.06p PD=615.6u AS=996.9525p PS=691.2u 
* M34 DRAIN GATE SOURCE BULK (257 14 259 88.5) 
M35 OUT IN VDD VDD CMOSP L=0.6u W=22.35u AD=885.06p PD=615.6u AS=996.9525p PS=691.2u 
* M35 DRAIN GATE SOURCE BULK (244 14 246 88.5) 
M36 OUT IN VDD VDD CMOSP L=0.6u W=22.35u AD=885.06p PD=615.6u AS=996.9525p PS=691.2u 
* M36 DRAIN GATE SOURCE BULK (231 14 233 88.5) 
M37 OUT IN VDD VDD CMOSP L=0.6u W=22.35u AD=885.06p PD=615.6u AS=996.9525p PS=691.2u 
* M37 DRAIN GATE SOURCE BULK (218 14 220 88.5) 
M38 OUT IN VDD VDD CMOSP L=0.6u W=22.35u AD=885.06p PD=615.6u AS=996.9525p PS=691.2u 
* M38 DRAIN GATE SOURCE BULK (205 14 207 88.5) 
M39 OUT IN VDD VDD CMOSP L=0.6u W=22.35u AD=885.06p PD=615.6u AS=996.9525p PS=691.2u 
* M39 DRAIN GATE SOURCE BULK (192 14 194 88.5) 
M40 OUT IN VDD VDD CMOSP L=0.6u W=22.35u AD=885.06p PD=615.6u AS=996.9525p PS=691.2u 
* M40 DRAIN GATE SOURCE BULK (179 14 181 88.5) 
M41 OUT IN VDD VDD CMOSP L=0.6u W=22.35u AD=885.06p PD=615.6u AS=996.9525p PS=691.2u 
* M41 DRAIN GATE SOURCE BULK (166 14 168 88.5) 
M42 OUT IN VDD VDD CMOSP L=0.6u W=22.35u AD=885.06p PD=615.6u AS=996.9525p PS=691.2u 
* M42 DRAIN GATE SOURCE BULK (153 14 155 88.5) 
M43 OUT IN VDD VDD CMOSP L=0.6u W=22.35u AD=885.06p PD=615.6u AS=996.9525p PS=691.2u 
* M43 DRAIN GATE SOURCE BULK (140 14 142 88.5) 
M44 OUT IN VDD VDD CMOSP L=0.6u W=22.35u AD=885.06p PD=615.6u AS=996.9525p PS=691.2u 
* M44 DRAIN GATE SOURCE BULK (127 14 129 88.5) 
M45 OUT IN VDD VDD CMOSP L=0.6u W=22.35u AD=885.06p PD=615.6u AS=996.9525p PS=691.2u 
* M45 DRAIN GATE SOURCE BULK (114 14 116 88.5) 
M46 OUT IN VDD VDD CMOSP L=0.6u W=22.35u AD=885.06p PD=615.6u AS=996.9525p PS=691.2u 
* M46 DRAIN GATE SOURCE BULK (101 14 103 88.5) 
M47 OUT IN VDD VDD CMOSP L=0.6u W=22.35u AD=885.06p PD=615.6u AS=996.9525p PS=691.2u 
* M47 DRAIN GATE SOURCE BULK (88 14 90 88.5) 
M48 OUT IN VDD VDD CMOSP L=0.6u W=22.35u AD=885.06p PD=615.6u AS=996.9525p PS=691.2u 
* M48 DRAIN GATE SOURCE BULK (75 14 77 88.5) 
M49 OUT IN VDD VDD CMOSP L=0.6u W=22.35u AD=885.06p PD=615.6u AS=996.9525p PS=691.2u 
* M49 DRAIN GATE SOURCE BULK (62 14 64 88.5) 
M50 OUT IN VDD VDD CMOSP L=0.6u W=22.35u AD=885.06p PD=615.6u AS=996.9525p PS=691.2u 
* M50 DRAIN GATE SOURCE BULK (49 14 51 88.5) 
M51 OUT IN VDD VDD CMOSP L=0.6u W=22.35u AD=885.06p PD=615.6u AS=996.9525p PS=691.2u 
* M51 DRAIN GATE SOURCE BULK (36 14 38 88.5) 
M52 OUT IN VDD VDD CMOSP L=0.6u W=22.35u AD=885.06p PD=615.6u AS=996.9525p PS=691.2u 
* M52 DRAIN GATE SOURCE BULK (23 14 25 88.5) 

* Total Nodes: 4
* Total Elements: 52
* Extract Elapsed Time: 2 seconds
.ENDS
