.SUBCKT INV IN OUT VDD GND
.param X=1 * X is drive strength(width multiplier), as in INVX1, INVX4, etc.

* OUT = ~IN

Mp OUT IN VDD VDD CMOSP
+L=0.6u 
+W=X*BALANCED_RATIO*MIN_CHANNEL_WIDTH
+AS=X*BALANCED_RATIO*MIN_CHANNEL_WIDTH*1.5u
+AD=X*BALANCED_RATIO*MIN_CHANNEL_WIDTH*1.5u
+PS=2.4u+(X*BALANCED_RATIO*MIN_CHANNEL_WIDTH*2)
+PD=2.4u+(X*BALANCED_RATIO*MIN_CHANNEL_WIDTH*2)

Mn OUT IN GND GND CMOSN 
+L=0.6u
+W=X*MIN_CHANNEL_WIDTH
+AS=X*MIN_CHANNEL_WIDTH*1.5u
+AD=X*MIN_CHANNEL_WIDTH*1.5u
+PS=2.4u+(X*MIN_CHANNEL_WIDTH*2)
+PD=2.4u+(X*MIN_CHANNEL_WIDTH*2)

.ENDS