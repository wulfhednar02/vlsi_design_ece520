.SUBCKT 2TMUX P_IN N_IN SEL OUT

* if (sel==0) out=P_IN
* else out=N_IN

Mp P_IN SEL OUT Vdd CMOSP L=0.6u W={{MIN_CHANNEL_WIDTH * BALANCED_RATIO}}
Mn N_IN SEL OUT GND CMOSN L=0.6u W={{MIN_CHANNEL_WIDTH}}
.ENDS
